module fibonacci 
(
    // Declaração das portas
    //------------
    input reset, clock, f_en;
    output f_valid;
    output [15,0] f_out;
    //------------
);

endmodule